** sch_path: /home/subhransu/gitRepo/test/runs/RUN_2025-12-21_23-08-25/parameters/transient_response/run_2/tran.sch
**.subckt tran
V1 VSS GND 0
V2 VDD GND 1.8
V3 vin GND CACE{vin}
x1 VDD Vout vin VSS inverter
C1 Vout GND 1e-12 m=1
**** begin user architecture code



.control
tran 0.1n 5.000000000000001e-07
set wr_singlescale
wrdata /home/subhransu/gitRepo/test/runs/RUN_2025-12-21_23-08-25/parameters/transient_response/run_2/tran_2.data V(Vout) V(Vin)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/subhransu/gitRepo/test/xschem/inverter.sym # of pins=4
** sym_path: /home/subhransu/gitRepo/test/xschem/inverter.sym
** sch_path: /home/subhransu/gitRepo/test/xschem/inverter.sch
.subckt inverter VDD vo vin VSS
*.opin vo
*.iopin VDD
*.iopin VSS
*.ipin vin
XM3 vo vin VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 vo vin VDD VDD pfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
