** sch_path: /home/subhransu/gitRepo/test/runs/RUN_2025-12-08_21-02-35/parameters/dc_params/run_0/tran.sch
**.subckt tran
V1 VSS GND 0
V2 VDD GND CACE{vdd}
V3 vin GND 0 PULSE(0 3.3 0 1n 1n 10n 20n)
x1 net1 net2 net3 net4 inverter
**** begin user architecture code



.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice tt

.include /home/subhransu/gitRepo/test/netlist/schematic/inverter.spice

.temp -40

.option warn=1






.control

.tran 0.1n 50n

.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/subhransu/gitRepo/test/xschem/inverter.sym # of pins=4
** sym_path: /home/subhransu/gitRepo/test/xschem/inverter.sym
** sch_path: /home/subhransu/gitRepo/test/xschem/inverter.sch
.subckt inverter VDD vo vin VSS
*.opin vo
*.iopin VDD
*.iopin VSS
*.ipin vin
XM3 vo vin VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 vo vin VDD VDD pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
